----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/04/2019 02:06:42 PM
-- Design Name: 
-- Module Name: problem2 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity problem2 is
  Port (A_1, A_2, B_1, B_2, D_1 :   in std_logic;
        E_out                   :   out std_logic);
end problem2;

architecture Behavioral of problem2 is
begin
    process(A_1, A_2, B_1, B_2, D_1) is
    begin
        if (A_1='1' and A_2='1') or (B_1='1' or B_2='1') or (B_2='1' and not(D_1)='1') then
            E_out <= '1';
        else
            E_out <= '0';
        end if;
    end process;
end Behavioral;
